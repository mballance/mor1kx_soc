
`include "uvm_macros.svh"

package mor1kx_soc_alt_uvm_env_pkg;
	import uvm_pkg::*;

	`include "mor1kx_soc_alt_uvm_env.svh"
	
endpackage
