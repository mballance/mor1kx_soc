
package my_pkg;
  typedef struct packed {logic a; logic b} my_struct_t;

endpackage

