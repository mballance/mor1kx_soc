/****************************************************************************
 * mor1kx_cluster.sv
 ****************************************************************************/

/**
 * Module: mor1kx_cluster
 * 
 * TODO: Add module documentation
 */
module mor1kx_cluster #(
			parameter int				N_CORES=2
		) (
		);
	


endmodule


