

`include "uvm_macros.svh"
package mor1kx_uvm_tests_pkg;
	import uvm_pkg::*;
	import mor1kx_uvm_env_pkg::*;
	
	`include "mor1kx_uvm_test_base.svh"
	
endpackage
