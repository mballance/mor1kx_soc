
`include "uvm_macros.svh"

package mor1kx_uvm_env_pkg;
	import uvm_pkg::*;
//	import generic_sram_byte_en_agent_pkg::*;
//	import generic_rom_agent_pkg::*;
	import uart_serial_agent_pkg::*;
//	import uvm_sdv_pkg::*;
//	import uvm_sdv_dpi_pkg::*;
//	import types_pkg::*;
	import vmon_client_pkg::*;

//	`include "simple_dpi_sdv_connector.svh"
	`include "mor1kx_uvm_env.svh"
	
endpackage
