

`include "uvm_macros.svh"
package mor1kx_soc_gate_uvm_tests_pkg;
	import uvm_pkg::*;
	import mor1kx_soc_gate_uvm_env_pkg::*;
	
	`include "mor1kx_soc_gate_uvm_test_base.svh"
	
endpackage
